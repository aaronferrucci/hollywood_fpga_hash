
`timescale 1ns/1ns
`default_nettype none

module sim_top;
  test_pw_gen_tb tb();
  test_program pgm();
endmodule

`default_nettype wire

